//////////////////////slv_error_write
class write_err_seq extends uvm_sequence#(transaction);
  `uvm_object_utils(write_err_seq)
  
  transaction tr;
 
  function new(string name = "write_err_seq");
    super.new(name);
  endfunction
  
  virtual task body();
    repeat(300)
      begin
        tr = transaction::type_id::create("tr");
        tr.addr_c.constraint_mode(0);
        tr.addr_c_err.constraint_mode(1);
        
        start_item(tr);
        assert(tr.randomize() with {
            op == writed;
        });
        finish_item(tr);   
      end
  endtask
  
 
endclass