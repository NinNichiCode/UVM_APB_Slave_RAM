
class wr_bulk_rd_bulk_test extends base_test;
    `uvm_component_utils(wr_bulk_rd_bulk_test)
 
function new(input string inst = "wr_bulk_rd_bulk_test", uvm_component c);
    super.new(inst,c);
endfunction

wr_bulk_rd_bulk_seq seq; 
  
 
virtual task run_test_seq();
   seq   = wr_bulk_rd_bulk_seq::type_id::create("seq");
    seq.start(env.a.seqr);
endtask
endclass
 